module muxAluSrc1(
	
);
endmodule
